module main

fn main() {
	x := u16(5)
	println(x)
}
